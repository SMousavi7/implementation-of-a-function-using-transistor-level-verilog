include"function";

module func_tb();

	reg a, b, c, d, _a, _b, _c, _d;
	wire output1;
	func func(output1, a, b, c, d, _a, _b, _c, _d);

	initial begin
		a = 0; 
		b = 0; 
 		c = 0; 
		d = 0; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;
		#20;
		a = 0; 
		b = 0; 
 		c = 0; 
		d = 1; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;
		#20;
		a = 0; 
		b = 0; 
 		c = 1; 
		d = 0; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;
		#20;
		a = 0; 
		b = 0; 
 		c = 1; 
		d = 1; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;
		#20;
		a = 0; 
		b = 1; 
 		c = 0; 
		d = 0; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;
		#20;
		a = 0; 
		b = 1; 
 		c = 0; 
		d = 1; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;
		#20;
		a = 0; 
		b = 1; 
 		c = 1; 
		d = 0; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;
		#20;
		a = 0; 
		b = 1; 
 		c = 1; 
		d = 1; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;

		#20;
		a = 1; 
		b = 0; 
 		c = 0;
		d = 0; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;

		#20;
		a = 1; 
		b = 0; 
 		c = 0; 
		d = 1; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;

		#20;
		a = 1; 
		b = 0; 
 		c = 1; 
		d = 0; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;

		#20;
		a = 1; 
		b = 0; 
 		c = 1; 
		d = 1; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;

		#20;
		a = 1; 
		b = 1; 
 		c = 0; 
		d = 0; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;

		#20;
		a = 1; 
		b = 1; 
 		c = 0; 
		d = 1; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;

		#20;
		a = 1; 
		b = 1; 
 		c = 1; 
		d = 0; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;

		#20;
		a = 1; 
		b = 1; 
 		c = 1; 
		d = 1; 
		_a = ~a;
		_b = ~b;
		_c = ~c;
		_d = ~d;

		#20;
	end
endmodule
